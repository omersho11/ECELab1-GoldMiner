module MainMenuBitmap (
	input logic clk,
	input logic resetN,
	input logic [10:0] offsetX,
	input logic [10:0] offsetY,
	input logic enable,

	output logic drawingRequest,
	output logic [7:0] RGBout
);

localparam int OBJECT_NUMBER_OF_X_BITS = 7;
localparam int OBJECT_NUMBER_OF_Y_BITS = 6;

localparam int OBJECT_HEIGHT_Y = 1 << OBJECT_NUMBER_OF_Y_BITS;
localparam int OBJECT_WIDTH_X  = 1 << OBJECT_NUMBER_OF_X_BITS;

logic [0:OBJECT_HEIGHT_Y-1][0:OBJECT_WIDTH_X-1][7:0] mainMenuColors = {

	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hfc, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd1, 8'hd5, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hf4, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hf8, 8'hfc, 8'hfc, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd0, 8'hd0, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd4, 8'hd4, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hf8, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd0, 8'hfc, 8'hf8, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfd, 8'hfd, 8'hd0, 8'hd0, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd0, 8'hd0, 8'hfd, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hf4, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd4, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hd1, 8'hf5, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hd1, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hf5, 8'hd5, 8'hd1, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc},
	{8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc, 8'hfc}
};







always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;
	end
	else begin
	if (enable) begin	
			drawingRequest <= 1'b1;
			RGBout <= (mainMenuColors[offsetY][offsetX]); 
		end
	end 
end

endmodule