module RotationTable #( 
	COUNT_SIZE = 8  // size of the table (in bits) 
)	
(	
	input	logic [COUNT_SIZE-1:0]	angle,
	
	output logic [7:0] sin,
	output logic sinIsNegative,
	output logic [7:0] cos,
	output logic cosIsNegative
);

localparam int table_size = (2**COUNT_SIZE)-1;
localparam int HALF_PI = 64;
localparam int PI = 128;
localparam int THREE_HALF_PI = 192;

logic [COUNT_SIZE-1:0] cosAngle;
assign cosAngle = angle + HALF_PI;

const logic [0:table_size-1] [7:0] sinTable = {
8'h0,
8'h6,
8'hC,
8'h12,
8'h18,
8'h1F,
8'h25,
8'h2B,
8'h31,
8'h37,
8'h3D,
8'h44,
8'h4A,
8'h4F,
8'h55,
8'h5B,
8'h61,
8'h67,
8'h6D,
8'h72,
8'h78,
8'h7D,
8'h83,
8'h88,
8'h8D,
8'h92,
8'h97,
8'h9C,
8'hA1,
8'hA6,
8'hAB,
8'hAF,
8'hB4,
8'hB8,
8'hBC,
8'hC1,
8'hC5,
8'hC9,
8'hCC,
8'hD0,
8'hD4,
8'hD7,
8'hDA,
8'hDD,
8'hE0,
8'hE3,
8'hE6,
8'hE9,
8'hEB,
8'hED,
8'hF0,
8'hF2,
8'hF4,
8'hF5,
8'hF7,
8'hF8,
8'hFA,
8'hFB,
8'hFC,
8'hFD,
8'hFD,
8'hFE,
8'hFE,
8'hFE,
8'hFF,
8'hFE,
8'hFE,
8'hFE,
8'hFD,
8'hFD,
8'hFC,
8'hFB,
8'hFA,
8'hF8,
8'hF7,
8'hF5,
8'hF4,
8'hF2,
8'hF0,
8'hED,
8'hEB,
8'hE9,
8'hE6,
8'hE3,
8'hE0,
8'hDD,
8'hDA,
8'hD7,
8'hD4,
8'hD0,
8'hCC,
8'hC9,
8'hC5,
8'hC1,
8'hBC,
8'hB8,
8'hB4,
8'hAF,
8'hAB,
8'hA6,
8'hA1,
8'h9C,
8'h97,
8'h92,
8'h8D,
8'h88,
8'h83,
8'h7D,
8'h78,
8'h72,
8'h6D,
8'h67,
8'h61,
8'h5B,
8'h55,
8'h4F,
8'h4A,
8'h44,
8'h3D,
8'h37,
8'h31,
8'h2B,
8'h25,
8'h1F,
8'h18,
8'h12,
8'hC,
8'h6,
8'h0,
8'h6,
8'hC,
8'h12,
8'h18,
8'h1F,
8'h25,
8'h2B,
8'h31,
8'h37,
8'h3D,
8'h44,
8'h4A,
8'h4F,
8'h55,
8'h5B,
8'h61,
8'h67,
8'h6D,
8'h72,
8'h78,
8'h7D,
8'h83,
8'h88,
8'h8D,
8'h92,
8'h97,
8'h9C,
8'hA1,
8'hA6,
8'hAB,
8'hAF,
8'hB4,
8'hB8,
8'hBC,
8'hC1,
8'hC5,
8'hC9,
8'hCC,
8'hD0,
8'hD4,
8'hD7,
8'hDA,
8'hDD,
8'hE0,
8'hE3,
8'hE6,
8'hE9,
8'hEB,
8'hED,
8'hF0,
8'hF2,
8'hF4,
8'hF5,
8'hF7,
8'hF8,
8'hFA,
8'hFB,
8'hFC,
8'hFD,
8'hFD,
8'hFE,
8'hFE,
8'hFE,
8'hFF,
8'hFE,
8'hFE,
8'hFE,
8'hFD,
8'hFD,
8'hFC,
8'hFB,
8'hFA,
8'hF8,
8'hF7,
8'hF5,
8'hF4,
8'hF2,
8'hF0,
8'hED,
8'hEB,
8'hE9,
8'hE6,
8'hE3,
8'hE0,
8'hDD,
8'hDA,
8'hD7,
8'hD4,
8'hD0,
8'hCC,
8'hC9,
8'hC5,
8'hC1,
8'hBC,
8'hB8,
8'hB4,
8'hAF,
8'hAB,
8'hA6,
8'hA1,
8'h9C,
8'h97,
8'h92,
8'h8D,
8'h88,
8'h83,
8'h7D,
8'h78,
8'h72,
8'h6D,
8'h67,
8'h61,
8'h5B,
8'h55,
8'h4F,
8'h4A,
8'h44,
8'h3D,
8'h37,
8'h31,
8'h2B,
8'h25,
8'h1F,
8'h18,
8'h12,
8'hC,
8'h6
};
 
//

always_comb begin

    // Shift the 8-bit signed value up to the top of the 16-bit signal
    sin = sinTable[angle]; 
    cos = sinTable[cosAngle];
	 sinIsNegative = angle > PI;
	 cosIsNegative = cosAngle > PI;
	 
end

endmodule